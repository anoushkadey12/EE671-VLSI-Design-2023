Question 1
.include models-180nm
*Name: Anoushka Dey
*Roll no: 210010010 :  nn = 10

*Rise and Fall times to achieve: 200+2*10=220 ps

*Parameters
*geometry parameters
.param pw = 1.865U
.param pl = 0.18U
.param pad = {2*pw*pl}
.param pas = {2*pw*pl}
.param ppd = {2*(pw + 2*pl)}
.param pps = {2*(pw + 2*pl)}

.param nw = 0.6465U
.param nl = 0.18U
.param nad = {2*nw*nl}
.param nas = {2*nw*nl}
.param npd = {2*(nw + 2*nl)}
.param nps = {2*(nw + 2*nl)}

* Minimum Inverter
.subckt inv supply Inp Output
*  This subcircuit defines a CMOS inverter with equal n and p widths
MP1 Output Inp Supply Supply cmosp
+ L={pl} W={pw} AD={pad} AS={pas} PD={ppd} PS={pps}
MN1 Output Inp 0      0      cmosn
+ L={nl} W={nw} AD={nad} AS={nas} PD={npd} PS={nps}
.ends

vdd supply 0 dc 1.8

*  Device under test
x3  supply Ck dutout inv

* Load Capacitor
C3 dutout 0 0.05pF


*TRANSIENT ANALYSIS with pulse inputs
VCk  Ck   0 DC 0 PULSE(0 1.8 0nS 20pS 20pS 4nS 8.0nS)
.tran 1pS 35nS 0nS

.control
run
plot 4.0+V(Ck) V(dutout)
meas tran inrise TRIG v(ck) VAL=0.18 RISE=2 TARG v(Ck) VAL=1.62 RISE=2
meas tran infall TRIG v(ck) VAL=1.62 FALL=2 TARG v(Ck) VAL=0.18 FALL=2
meas tran drise TRIG v(dutout) VAL=0.18 RISE=2 TARG v(dutout) VAL=1.62 RISE=2
meas tran dfall TRIG v(dutout) VAL=1.62 FALL=2 TARG v(dutout) VAL=0.18 FALL=2
.endc
.end
