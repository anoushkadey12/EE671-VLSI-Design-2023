Assignment 2
.include models-180nm
*Name: Anoushka Dey
*Roll 210010010 :  nn = 10

*Rise and Fall times to achieve: 200+2*10=220 ps

*Parameters
*geometry parameters
.param pw = 1.865U
.param pl = 0.18U
.param pad = {2*pw*pl}
.param pas = {2*pw*pl}
.param ppd = {2*(pw + 2*pl)}
.param pps = {2*(pw + 2*pl)}

.param nw = 0.6465U
.param nl = 0.18U
.param nad = {2*nw*nl}
.param nas = {2*nw*nl}
.param npd = {2*(nw + 2*nl)}
.param nps = {2*(nw + 2*nl)}

* Minimum Inverter
.subckt inv supply Inp Output
*  This subcircuit defines a CMOS inverter with equal n and p widths
MP1 Output Inp Supply Supply cmosp
+ L={pl} W={pw} AD={pad} AS={pas} PD={ppd} PS={pps}
MN1 Output Inp 0      0      cmosn
+ L={nl} W={nw} AD={nad} AS={nas} PD={npd} PS={nps}
.ends

*Input Shaper
* pulse with time period of Trep, rise and fall times = Trep/20
.param Trep= 5n
.param Trf = {Trep/20.0}
.param Tw = {Trep/2.0 - Trf}
.param hival=1.8
.param loval=0.0
Vpulse pgen 0 DC 0 PULSE({loval} {hival} {Tw} {Trf} {Trf} {Tw} {Trep})


vdd supply 0 dc 1.8
xinvstart supply pgen node1 inv
xinv1 supply node1 node2 inv
xinv2 supply node2 dutin inv
xinv3 supply node2 node3 inv
xinv4 supply node2 node3 inv
xinv5 supply node2 node3 inv
C1 node3 0 0.1p

*Device Under Test
xdut supply dutin dutout inv

*Test Load
xinv6 supply dutout node5 inv
xinv7 supply dutout node5 inv
*xinv8 supply dutout node5 inv
*xinv9 supply dutout node5 inv
*xinv10 supply dutout node5 inv
*xinv11 supply dutout node5 inv
*xinv12 supply dutout node5 inv
*xinv13 supply dutout node5 inv

*Load on load
xinv14 supply node5 node6 inv
xinv15 supply node5 node6 inv
xinv16 supply node5 node6 inv
xinv17 supply node5 node6 inv
C2 node6 0 0.1p

.tran 1pS {3*Trep} 0nS
.control
run
meas tran rise_delay TRIG v(dutin) VAL=0.9 RISE=2 TARG v(dutout) VAL=0.9 FALL=2
meas tran fall_delay TRIG v(dutin) VAL=0.9 FALL=2 TARG v(dutout) VAL=0.9 RISE=2
let delay={(rise_delay+fall_delay)/2}
print delay
.endc
.end



